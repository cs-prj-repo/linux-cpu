module execute(

);


endmodule