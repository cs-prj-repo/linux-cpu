module reg_if1_if2(
    

);


endmodule