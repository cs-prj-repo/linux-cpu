module satp(

);
reg [63:0] satp;
reg [63:0] 

always 

reg [63:0] mcpuid;
reg [63:0] mimpid;
reg [63:0] mhartid;
reg [63:0] mstatus;
reg [63:0] mtvex;
reg [63:0] mtdeleg;
reg [63:0] mip;
reg [63:0] mie;
reg [63:0] mtime;
reg [63:0] mtimecmp;
reg [63:0] mscratch;
reg [63:0] mepc;
reg [63:0] mcause;
reg [63:0] mbadaddr;
reg [63:0] sstatus;

endmodule