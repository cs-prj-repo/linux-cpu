module regW(
    input wire memory_i_mem_data;
);


endmodule