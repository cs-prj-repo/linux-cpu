module regE(
    input  wire clk,
    input  wire rst,
    input  wire decode_i_bus_info,
    output wire regE_o_bus_info
);
always @(posedge clk) begin
    if(rst) begin
        
    end
    else begin
 
    end
end
endmodule