module execute(
    input  wire [63:0] regD_i_regdata1,
    input  wire [63:0] regD_i_regdata2,
    output wire [63:0] execute_o_alu_result
);


endmodule