module regW(
    input wire clk,
    input wire rst,
    input wire regM_i_bus_info,
    input wire regM_i_commit_info,
    output reg regW_o_bus_info,
    output reg regW_o_commit_info
);
always @(posedge clk) begin
    if(rst) begin
        
    end
    else begin
        
    end
end

endmodule