module decode(
    input wire regD_i_bus_info
);


endmodule