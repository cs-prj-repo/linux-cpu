module decode(
    input  wire [95:0] regD_i_bus_info,
    output wire decode_o_bus_info
);


endmodule