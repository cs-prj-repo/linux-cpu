module regE(
    input wire decode_i_
    input wire decode_


);

endmodule