module execute(
    input  wire regE_i_bus_info,
    input  wire regE_i_commit_info,

    output wire execute_o_bus_info,
    output wire execute_o_commit_info
);


endmodule