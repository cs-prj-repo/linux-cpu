module write_back(
    input wire regW_i_bus_info
);


endmodule