module fetch(
    input  wire   pc_o_bus,
    output wire   fetch_o_bus
);


endmodule